module naive (
    input A, B, C, D,
    output Y
);

assign Y = ; // Enter your equation here

endmodule
